module example (a, b, c, y);
  input a;
  input b;
  input c;  
  output y;
endmodule

/* 
* A module is the main building block in Verilog
*
* So, what we need to declare it?
* Just:
* - Name of the module
* - Types of its connections (input, output)
* - Name of its connection
* */
